module Data_Hazard_Detect();

// Assuming we have X to X forwarding, the only data hazard
// we need to watch out for is RAW, Branching


endmodule