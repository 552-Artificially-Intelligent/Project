module M_W_Flops();




endmodule