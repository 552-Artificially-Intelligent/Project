module D_X_Flops(clk, rst, en,
		oldPC_in, new_PC_in, oldPC_out, new_PC_out,
		
		);





endmodule