module M_W_Flops(clk, rst, en,);

input clk, rst, en, 

// Data


// Signals


endmodule