module Data_Hazard_Detect();




endmodule