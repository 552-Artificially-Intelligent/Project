module D_X_Flops(clk, rst, en,
		,

		);





endmodule