module Forwarding_Unit(
	X_M_RegWrite, X_M_MemWrite,
	M_W_RegWrite, 



);






endmodule