module D_X_Flops(
	clk, rst, en,
	// Signals
	D_ALUsrc, D_X_ALUsrc,
	D_MemtoReg, D_X_MemtoReg,
	D_RegWrite, D_X_RegWrite,
	D_MemRead, D_X_MemRead,
	D_MemWrite, D_X_MemWrite,
	D_branch_inst, D_X_branch_inst,
	D_branch_src, D_X_branch_src,
	D_RegDst, D_X_RegDst,
	D_SavePC, D_X_SavePC,
	F_D_halt, D_X_halt,

	// Data
	

);
// TODO





endmodule