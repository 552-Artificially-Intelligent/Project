module X_M_Flops();





endmodule